library verilog;
use verilog.vl_types.all;
entity Projeto3U_vlg_vec_tst is
end Projeto3U_vlg_vec_tst;
