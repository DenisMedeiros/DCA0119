library verilog;
use verilog.vl_types.all;
entity Projeto3U_vlg_sample_tst is
    port(
        CLOCK_50MHZ     : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Projeto3U_vlg_sample_tst;
