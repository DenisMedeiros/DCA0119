library verilog;
use verilog.vl_types.all;
entity Projeto3U_vlg_check_tst is
    port(
        CLOCK_50KHZ     : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Projeto3U_vlg_check_tst;
