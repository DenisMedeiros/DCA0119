library verilog;
use verilog.vl_types.all;
entity Projeto3U is
    port(
        CLOCK_50KHZ     : out    vl_logic;
        CLOCK_50MHZ     : in     vl_logic
    );
end Projeto3U;
